/////////////////////////////////////////////////
// ��ģ��
/////////////////////////////////////////////////

module led(
    input       clk,
    input       rst,
    input       
);