#
# ��֤ƽ̨����
#

module partfreq_test(
    input       clk,
    input       rst,
    output      clk_out
);

    .clk        (clk),
    .rst        (rst),
    .clk_out    (clk_out)