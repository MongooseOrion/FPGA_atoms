//
// UART ����ģ��
//
//
module uart_trans #(
    parameter UART_BOT = 'd9600
)(
    input           sys_clk,
    input           sys_rst
);


endmodule