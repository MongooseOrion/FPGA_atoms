//
// SDRAM ������ģ��
/* SDRAMҳͻ���������ľ������̣�
1. ���ͼ���ָ�SDRAM��ͬʱBA0-BA1��A0-A12�ֱ�д��L-Bank��ַ���е�ַ�������ض�L-Bank���ض��У�
2. ����ָ��д��󣬵ȴ�tRCDʱ�䣬�˹����в��������Ϊ�ղ������
3. tRCD�ȴ�ʱ�������д�������ָ�ͬʱA0-A8д�����ݶ�ȡ�׵�ַ��
4. ������ָ��д��������ת��Ǳ��״̬���ȴ�Ǳ���ڽ�����DQ��ʼ�����ȡ���ݣ����ȡ���ݸ���ΪN��
5. �Զ�ָ��д�����ڵ��¸�ʱ�����ڿ�ʼ������N��ʱ�����ں�д��ͻ��ָֹͣ���ֹ���ݶ�������
6. ͻ��ָֹͣ��д���DQ������������������ɺ�SDRAM��ҳͻ����������ɡ�
*/
//

module sdram_read(
    input               sys_clk,
    input               sys_rst,
    input               init_end,
    input               rd_en,
    input      [23:0]   rd_addr,
    input      [15:0]   rd_data,

    output              rd_ack,
    output              rd_end,
    output reg []
);