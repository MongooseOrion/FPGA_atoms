module muxtwo(
    
)