//
// SDRAM ��ʼ��ģ��
/* SDRAM ��ʼ�����̣�
    1. �� SDRAM �ϵ磬�����ȶ�ʱ���źţ�CKE ����Ϊ�ߵ�ƽ��
    2. �ȴ� T>=100us ��ʱ�䣬�˹����в��������Ϊ�ղ������
    3. 100us�ȴ�������д��Ԥ������A10����Ϊ�ߵ�ƽ��������L-Bank����Ԥ��磻
    4. Ԥ���ָ��д��󣬵ȴ�tRPʱ�䣬�˹����в��������Ϊ�ղ������
    5. tRP�ȴ�ʱ�������д���Զ�ˢ�����
    6. �Զ�ˢ������д��󣬵ȴ�tRCʱ�䣬�˹����в��������Ϊ�ղ������
    7. tRC�ȴ�ʱ��������ٴ�д���Զ�ˢ�����
    8. �Զ�ˢ������д��󣬵ȴ�tRCʱ�䣬�˹����в��������Ϊ�ղ������
    9. tRC�ȴ�ʱ�������д��ģʽ�Ĵ�������ָ���ַ����A0-A11������ͬ����ģʽ�Ĵ�����ͬģʽ�����ã�
    10. ģʽ�Ĵ�������ָ��д��󣬵ȴ�tMRDʱ�䣬�˹����в��������Ϊ�ղ������
    11. tMRD�ȴ�ʱ�������SDRAM��ʼ����ɡ�
*/
//
//

module sdram_init #()(

    input               sys_clk,    // 100MHz
    input               sys_rst,

    output reg [3:0]    init_cmd,
    output reg [1:0]    init_ba,
    output reg [12:0]   init_addr,
    output              init_end
);

localparam  T_POWER = 15'd20_000;   // �����ϵ�ʱ�ӵȴ� 200us
localparam  P_CHARGE = 4'b0010,     // Ԥ���ָ��
            AUTO_REF = 4'b0001,     // �Զ�ˢ��ָ��
            NOP = 4'b0111 ,         // �ղ���ָ��
            M_REG_SET = 4'b0000 ;   // ģʽ�Ĵ�������ָ��

// SDRAM��ʼ�����̸���״̬
localparam  INIT_IDLE = 3'b000 ,    //��ʼ״̬
            INIT_PRE = 3'b001 ,     //Ԥ���״̬
            INIT_TRP = 3'b011 ,     //Ԥ���ȴ� tRP
            INIT_AR = 3'b010 ,      //�Զ�ˢ��
            INIT_TRF = 3'b100 ,     //�Զ�ˢ�µȴ� tRC
            INIT_MRS = 3'b101 ,     //ģʽ�Ĵ�������
            INIT_TMRD = 3'b111 ,    //ģʽ�Ĵ������õȴ� tMRD
            INIT_END = 3'b110 ;     //��ʼ�����

localparam  TRP_CLK = 3'd2 ,        //Ԥ���ȴ�����,20ns
            TRC_CLK = 3'd7 ,        //�Զ�ˢ�µȴ�,70ns
            TMRD_CLK = 3'd3 ;       //ģʽ�Ĵ������õȴ�����,30ns

reg 